module Vector2(
  input  [31:0] io_in,
  output [31:0] io_out
);
  io_out_hi,io_out_lo}; // @[Cat.scala 30:58]
endmodule
