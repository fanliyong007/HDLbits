module Wire(
  input   in,
  output  out
);
  assign out = in; // @[Wire.scala 11:10]
endmodule
