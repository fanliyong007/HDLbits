module FullAdder(
  input   io_a,
  input   io_b,
  input   io_cin,
  output  io_sum,
  output  io_cout
);
  wire  a_xor_b = io_a ^ io_b; // @[FullAdder.scala 15:22]
  wire  a_and_b = io_a & io_b; // @[FullAdder.scala 18:22]
  wire  b_and_cin = io_b & io_cin; // @[FullAdder.scala 19:24]
  wire  a_and_cin = io_a & io_cin; // @[FullAdder.scala 20:24]
  assign io_sum = a_xor_b ^ io_cin; // @[FullAdder.scala 16:21]
  assign io_cout = a_and_b | b_and_cin | a_and_cin; // @[FullAdder.scala 21:34]
endmodule
module Adder(
  input  [99:0] io_A,
  input  [99:0] io_B,
  input         io_Cin,
  output [99:0] io_Sum,
  output [99:0] io_Cout
);
  wire  FullAdder_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_1_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_1_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_1_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_1_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_1_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_2_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_2_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_2_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_2_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_2_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_3_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_3_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_3_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_3_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_3_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_4_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_4_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_4_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_4_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_4_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_5_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_5_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_5_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_5_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_5_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_6_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_6_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_6_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_6_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_6_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_7_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_7_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_7_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_7_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_7_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_8_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_8_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_8_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_8_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_8_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_9_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_9_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_9_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_9_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_9_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_10_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_10_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_10_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_10_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_10_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_11_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_11_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_11_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_11_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_11_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_12_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_12_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_12_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_12_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_12_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_13_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_13_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_13_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_13_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_13_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_14_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_14_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_14_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_14_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_14_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_15_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_15_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_15_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_15_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_15_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_16_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_16_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_16_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_16_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_16_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_17_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_17_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_17_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_17_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_17_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_18_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_18_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_18_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_18_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_18_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_19_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_19_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_19_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_19_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_19_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_20_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_20_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_20_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_20_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_20_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_21_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_21_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_21_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_21_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_21_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_22_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_22_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_22_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_22_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_22_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_23_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_23_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_23_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_23_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_23_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_24_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_24_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_24_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_24_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_24_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_25_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_25_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_25_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_25_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_25_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_26_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_26_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_26_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_26_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_26_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_27_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_27_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_27_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_27_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_27_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_28_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_28_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_28_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_28_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_28_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_29_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_29_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_29_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_29_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_29_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_30_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_30_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_30_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_30_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_30_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_31_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_31_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_31_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_31_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_31_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_32_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_32_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_32_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_32_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_32_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_33_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_33_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_33_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_33_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_33_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_34_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_34_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_34_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_34_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_34_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_35_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_35_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_35_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_35_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_35_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_36_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_36_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_36_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_36_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_36_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_37_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_37_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_37_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_37_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_37_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_38_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_38_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_38_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_38_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_38_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_39_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_39_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_39_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_39_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_39_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_40_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_40_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_40_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_40_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_40_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_41_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_41_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_41_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_41_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_41_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_42_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_42_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_42_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_42_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_42_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_43_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_43_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_43_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_43_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_43_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_44_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_44_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_44_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_44_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_44_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_45_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_45_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_45_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_45_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_45_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_46_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_46_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_46_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_46_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_46_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_47_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_47_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_47_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_47_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_47_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_48_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_48_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_48_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_48_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_48_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_49_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_49_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_49_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_49_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_49_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_50_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_50_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_50_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_50_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_50_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_51_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_51_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_51_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_51_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_51_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_52_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_52_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_52_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_52_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_52_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_53_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_53_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_53_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_53_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_53_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_54_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_54_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_54_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_54_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_54_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_55_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_55_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_55_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_55_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_55_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_56_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_56_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_56_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_56_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_56_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_57_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_57_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_57_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_57_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_57_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_58_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_58_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_58_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_58_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_58_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_59_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_59_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_59_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_59_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_59_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_60_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_60_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_60_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_60_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_60_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_61_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_61_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_61_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_61_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_61_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_62_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_62_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_62_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_62_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_62_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_63_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_63_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_63_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_63_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_63_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_64_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_64_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_64_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_64_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_64_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_65_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_65_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_65_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_65_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_65_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_66_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_66_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_66_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_66_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_66_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_67_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_67_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_67_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_67_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_67_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_68_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_68_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_68_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_68_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_68_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_69_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_69_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_69_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_69_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_69_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_70_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_70_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_70_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_70_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_70_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_71_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_71_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_71_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_71_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_71_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_72_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_72_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_72_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_72_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_72_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_73_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_73_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_73_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_73_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_73_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_74_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_74_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_74_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_74_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_74_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_75_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_75_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_75_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_75_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_75_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_76_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_76_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_76_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_76_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_76_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_77_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_77_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_77_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_77_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_77_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_78_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_78_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_78_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_78_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_78_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_79_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_79_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_79_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_79_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_79_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_80_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_80_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_80_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_80_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_80_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_81_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_81_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_81_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_81_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_81_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_82_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_82_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_82_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_82_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_82_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_83_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_83_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_83_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_83_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_83_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_84_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_84_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_84_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_84_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_84_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_85_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_85_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_85_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_85_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_85_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_86_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_86_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_86_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_86_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_86_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_87_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_87_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_87_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_87_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_87_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_88_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_88_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_88_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_88_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_88_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_89_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_89_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_89_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_89_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_89_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_90_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_90_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_90_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_90_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_90_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_91_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_91_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_91_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_91_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_91_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_92_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_92_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_92_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_92_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_92_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_93_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_93_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_93_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_93_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_93_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_94_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_94_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_94_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_94_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_94_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_95_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_95_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_95_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_95_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_95_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_96_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_96_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_96_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_96_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_96_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_97_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_97_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_97_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_97_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_97_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_98_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_98_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_98_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_98_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_98_io_cout; // @[Adder.scala 19:35]
  wire  FullAdder_99_io_a; // @[Adder.scala 19:35]
  wire  FullAdder_99_io_b; // @[Adder.scala 19:35]
  wire  FullAdder_99_io_cin; // @[Adder.scala 19:35]
  wire  FullAdder_99_io_sum; // @[Adder.scala 19:35]
  wire  FullAdder_99_io_cout; // @[Adder.scala 19:35]
  wire  sum_0 = FullAdder_io_sum; // @[Adder.scala 32:26]
  wire  sum_1 = FullAdder_1_io_sum; // @[Adder.scala 32:26]
  wire  sum_2 = FullAdder_2_io_sum; // @[Adder.scala 32:26]
  wire  sum_3 = FullAdder_3_io_sum; // @[Adder.scala 32:26]
  wire  sum_4 = FullAdder_4_io_sum; // @[Adder.scala 32:26]
  wire  sum_5 = FullAdder_5_io_sum; // @[Adder.scala 32:26]
  wire  sum_6 = FullAdder_6_io_sum; // @[Adder.scala 32:26]
  wire  sum_7 = FullAdder_7_io_sum; // @[Adder.scala 32:26]
  wire  sum_8 = FullAdder_8_io_sum; // @[Adder.scala 32:26]
  wire  sum_9 = FullAdder_9_io_sum; // @[Adder.scala 32:26]
  wire  sum_10 = FullAdder_10_io_sum; // @[Adder.scala 32:26]
  wire  sum_11 = FullAdder_11_io_sum; // @[Adder.scala 32:26]
  wire  sum_12 = FullAdder_12_io_sum; // @[Adder.scala 32:26]
  wire  sum_13 = FullAdder_13_io_sum; // @[Adder.scala 32:26]
  wire  sum_14 = FullAdder_14_io_sum; // @[Adder.scala 32:26]
  wire  sum_15 = FullAdder_15_io_sum; // @[Adder.scala 32:26]
  wire  sum_16 = FullAdder_16_io_sum; // @[Adder.scala 32:26]
  wire  sum_17 = FullAdder_17_io_sum; // @[Adder.scala 32:26]
  wire  sum_18 = FullAdder_18_io_sum; // @[Adder.scala 32:26]
  wire  sum_19 = FullAdder_19_io_sum; // @[Adder.scala 32:26]
  wire  sum_20 = FullAdder_20_io_sum; // @[Adder.scala 32:26]
  wire  sum_21 = FullAdder_21_io_sum; // @[Adder.scala 32:26]
  wire  sum_22 = FullAdder_22_io_sum; // @[Adder.scala 32:26]
  wire  sum_23 = FullAdder_23_io_sum; // @[Adder.scala 32:26]
  wire  sum_24 = FullAdder_24_io_sum; // @[Adder.scala 32:26]
  wire  sum_25 = FullAdder_25_io_sum; // @[Adder.scala 32:26]
  wire  sum_26 = FullAdder_26_io_sum; // @[Adder.scala 32:26]
  wire  sum_27 = FullAdder_27_io_sum; // @[Adder.scala 32:26]
  wire  sum_28 = FullAdder_28_io_sum; // @[Adder.scala 32:26]
  wire  sum_29 = FullAdder_29_io_sum; // @[Adder.scala 32:26]
  wire  sum_30 = FullAdder_30_io_sum; // @[Adder.scala 32:26]
  wire  sum_31 = FullAdder_31_io_sum; // @[Adder.scala 32:26]
  wire  sum_32 = FullAdder_32_io_sum; // @[Adder.scala 32:26]
  wire  sum_33 = FullAdder_33_io_sum; // @[Adder.scala 32:26]
  wire  sum_34 = FullAdder_34_io_sum; // @[Adder.scala 32:26]
  wire  sum_35 = FullAdder_35_io_sum; // @[Adder.scala 32:26]
  wire  sum_36 = FullAdder_36_io_sum; // @[Adder.scala 32:26]
  wire  sum_37 = FullAdder_37_io_sum; // @[Adder.scala 32:26]
  wire  sum_38 = FullAdder_38_io_sum; // @[Adder.scala 32:26]
  wire  sum_39 = FullAdder_39_io_sum; // @[Adder.scala 32:26]
  wire  sum_40 = FullAdder_40_io_sum; // @[Adder.scala 32:26]
  wire  sum_41 = FullAdder_41_io_sum; // @[Adder.scala 32:26]
  wire  sum_42 = FullAdder_42_io_sum; // @[Adder.scala 32:26]
  wire  sum_43 = FullAdder_43_io_sum; // @[Adder.scala 32:26]
  wire  sum_44 = FullAdder_44_io_sum; // @[Adder.scala 32:26]
  wire  sum_45 = FullAdder_45_io_sum; // @[Adder.scala 32:26]
  wire  sum_46 = FullAdder_46_io_sum; // @[Adder.scala 32:26]
  wire  sum_47 = FullAdder_47_io_sum; // @[Adder.scala 32:26]
  wire  sum_48 = FullAdder_48_io_sum; // @[Adder.scala 32:26]
  wire  sum_49 = FullAdder_49_io_sum; // @[Adder.scala 32:26]
  wire  sum_50 = FullAdder_50_io_sum; // @[Adder.scala 32:26]
  wire  sum_51 = FullAdder_51_io_sum; // @[Adder.scala 32:26]
  wire  sum_52 = FullAdder_52_io_sum; // @[Adder.scala 32:26]
  wire  sum_53 = FullAdder_53_io_sum; // @[Adder.scala 32:26]
  wire  sum_54 = FullAdder_54_io_sum; // @[Adder.scala 32:26]
  wire  sum_55 = FullAdder_55_io_sum; // @[Adder.scala 32:26]
  wire  sum_56 = FullAdder_56_io_sum; // @[Adder.scala 32:26]
  wire  sum_57 = FullAdder_57_io_sum; // @[Adder.scala 32:26]
  wire  sum_58 = FullAdder_58_io_sum; // @[Adder.scala 32:26]
  wire  sum_59 = FullAdder_59_io_sum; // @[Adder.scala 32:26]
  wire  sum_60 = FullAdder_60_io_sum; // @[Adder.scala 32:26]
  wire  sum_61 = FullAdder_61_io_sum; // @[Adder.scala 32:26]
  wire  sum_62 = FullAdder_62_io_sum; // @[Adder.scala 32:26]
  wire  sum_63 = FullAdder_63_io_sum; // @[Adder.scala 32:26]
  wire  sum_64 = FullAdder_64_io_sum; // @[Adder.scala 32:26]
  wire  sum_65 = FullAdder_65_io_sum; // @[Adder.scala 32:26]
  wire  sum_66 = FullAdder_66_io_sum; // @[Adder.scala 32:26]
  wire  sum_67 = FullAdder_67_io_sum; // @[Adder.scala 32:26]
  wire  sum_68 = FullAdder_68_io_sum; // @[Adder.scala 32:26]
  wire  sum_69 = FullAdder_69_io_sum; // @[Adder.scala 32:26]
  wire  sum_70 = FullAdder_70_io_sum; // @[Adder.scala 32:26]
  wire  sum_71 = FullAdder_71_io_sum; // @[Adder.scala 32:26]
  wire  sum_72 = FullAdder_72_io_sum; // @[Adder.scala 32:26]
  wire  sum_73 = FullAdder_73_io_sum; // @[Adder.scala 32:26]
  wire  sum_74 = FullAdder_74_io_sum; // @[Adder.scala 32:26]
  wire  sum_75 = FullAdder_75_io_sum; // @[Adder.scala 32:26]
  wire  sum_76 = FullAdder_76_io_sum; // @[Adder.scala 32:26]
  wire  sum_77 = FullAdder_77_io_sum; // @[Adder.scala 32:26]
  wire  sum_78 = FullAdder_78_io_sum; // @[Adder.scala 32:26]
  wire  sum_79 = FullAdder_79_io_sum; // @[Adder.scala 32:26]
  wire  sum_80 = FullAdder_80_io_sum; // @[Adder.scala 32:26]
  wire  sum_81 = FullAdder_81_io_sum; // @[Adder.scala 32:26]
  wire  sum_82 = FullAdder_82_io_sum; // @[Adder.scala 32:26]
  wire  sum_83 = FullAdder_83_io_sum; // @[Adder.scala 32:26]
  wire  sum_84 = FullAdder_84_io_sum; // @[Adder.scala 32:26]
  wire  sum_85 = FullAdder_85_io_sum; // @[Adder.scala 32:26]
  wire  sum_86 = FullAdder_86_io_sum; // @[Adder.scala 32:26]
  wire  sum_87 = FullAdder_87_io_sum; // @[Adder.scala 32:26]
  wire  sum_88 = FullAdder_88_io_sum; // @[Adder.scala 32:26]
  wire  sum_89 = FullAdder_89_io_sum; // @[Adder.scala 32:26]
  wire  sum_90 = FullAdder_90_io_sum; // @[Adder.scala 32:26]
  wire  sum_91 = FullAdder_91_io_sum; // @[Adder.scala 32:26]
  wire  sum_92 = FullAdder_92_io_sum; // @[Adder.scala 32:26]
  wire  sum_93 = FullAdder_93_io_sum; // @[Adder.scala 32:26]
  wire  sum_94 = FullAdder_94_io_sum; // @[Adder.scala 32:26]
  wire  sum_95 = FullAdder_95_io_sum; // @[Adder.scala 32:26]
  wire  sum_96 = FullAdder_96_io_sum; // @[Adder.scala 32:26]
  wire  sum_97 = FullAdder_97_io_sum; // @[Adder.scala 32:26]
  wire  sum_98 = FullAdder_98_io_sum; // @[Adder.scala 32:26]
  wire  sum_99 = FullAdder_99_io_sum; // @[Adder.scala 32:26]
  wire [5:0] io_Sum_lo_lo_lo_lo = {sum_5,sum_4,sum_3,sum_2,sum_1,sum_0}; // @[Adder.scala 34:17]
  wire [11:0] io_Sum_lo_lo_lo = {sum_11,sum_10,sum_9,sum_8,sum_7,sum_6,io_Sum_lo_lo_lo_lo}; // @[Adder.scala 34:17]
  wire [5:0] io_Sum_lo_lo_hi_lo = {sum_17,sum_16,sum_15,sum_14,sum_13,sum_12}; // @[Adder.scala 34:17]
  wire [24:0] io_Sum_lo_lo = {sum_24,sum_23,sum_22,sum_21,sum_20,sum_19,sum_18,io_Sum_lo_lo_hi_lo,io_Sum_lo_lo_lo}; // @[Adder.scala 34:17]
  wire [5:0] io_Sum_lo_hi_lo_lo = {sum_30,sum_29,sum_28,sum_27,sum_26,sum_25}; // @[Adder.scala 34:17]
  wire [11:0] io_Sum_lo_hi_lo = {sum_36,sum_35,sum_34,sum_33,sum_32,sum_31,io_Sum_lo_hi_lo_lo}; // @[Adder.scala 34:17]
  wire [5:0] io_Sum_lo_hi_hi_lo = {sum_42,sum_41,sum_40,sum_39,sum_38,sum_37}; // @[Adder.scala 34:17]
  wire [49:0] io_Sum_lo = {sum_49,sum_48,sum_47,sum_46,sum_45,sum_44,sum_43,io_Sum_lo_hi_hi_lo,io_Sum_lo_hi_lo,
    io_Sum_lo_lo}; // @[Adder.scala 34:17]
  wire [5:0] io_Sum_hi_lo_lo_lo = {sum_55,sum_54,sum_53,sum_52,sum_51,sum_50}; // @[Adder.scala 34:17]
  wire [11:0] io_Sum_hi_lo_lo = {sum_61,sum_60,sum_59,sum_58,sum_57,sum_56,io_Sum_hi_lo_lo_lo}; // @[Adder.scala 34:17]
  wire [5:0] io_Sum_hi_lo_hi_lo = {sum_67,sum_66,sum_65,sum_64,sum_63,sum_62}; // @[Adder.scala 34:17]
  wire [24:0] io_Sum_hi_lo = {sum_74,sum_73,sum_72,sum_71,sum_70,sum_69,sum_68,io_Sum_hi_lo_hi_lo,io_Sum_hi_lo_lo}; // @[Adder.scala 34:17]
  wire [5:0] io_Sum_hi_hi_lo_lo = {sum_80,sum_79,sum_78,sum_77,sum_76,sum_75}; // @[Adder.scala 34:17]
  wire [11:0] io_Sum_hi_hi_lo = {sum_86,sum_85,sum_84,sum_83,sum_82,sum_81,io_Sum_hi_hi_lo_lo}; // @[Adder.scala 34:17]
  wire [5:0] io_Sum_hi_hi_hi_lo = {sum_92,sum_91,sum_90,sum_89,sum_88,sum_87}; // @[Adder.scala 34:17]
  wire [49:0] io_Sum_hi = {sum_99,sum_98,sum_97,sum_96,sum_95,sum_94,sum_93,io_Sum_hi_hi_hi_lo,io_Sum_hi_hi_lo,
    io_Sum_hi_lo}; // @[Adder.scala 34:17]
  wire  mycout_2 = FullAdder_2_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_1 = FullAdder_1_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_0 = FullAdder_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_5 = FullAdder_5_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_4 = FullAdder_4_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_3 = FullAdder_3_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_lo_lo_lo_lo = {mycout_5,mycout_4,mycout_3,mycout_2,mycout_1,mycout_0}; // @[Adder.scala 35:21]
  wire  mycout_8 = FullAdder_8_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_7 = FullAdder_7_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_6 = FullAdder_6_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_11 = FullAdder_11_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_10 = FullAdder_10_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_9 = FullAdder_9_io_cout; // @[Adder.scala 22:20 31:15]
  wire [11:0] io_Cout_lo_lo_lo = {mycout_11,mycout_10,mycout_9,mycout_8,mycout_7,mycout_6,io_Cout_lo_lo_lo_lo}; // @[Adder.scala 35:21]
  wire  mycout_14 = FullAdder_14_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_13 = FullAdder_13_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_12 = FullAdder_12_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_17 = FullAdder_17_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_16 = FullAdder_16_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_15 = FullAdder_15_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_lo_lo_hi_lo = {mycout_17,mycout_16,mycout_15,mycout_14,mycout_13,mycout_12}; // @[Adder.scala 35:21]
  wire  mycout_20 = FullAdder_20_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_19 = FullAdder_19_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_18 = FullAdder_18_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_22 = FullAdder_22_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_21 = FullAdder_21_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_24 = FullAdder_24_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_23 = FullAdder_23_io_cout; // @[Adder.scala 22:20 31:15]
  wire [24:0] io_Cout_lo_lo = {mycout_24,mycout_23,mycout_22,mycout_21,mycout_20,mycout_19,mycout_18,io_Cout_lo_lo_hi_lo
    ,io_Cout_lo_lo_lo}; // @[Adder.scala 35:21]
  wire  mycout_27 = FullAdder_27_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_26 = FullAdder_26_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_25 = FullAdder_25_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_30 = FullAdder_30_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_29 = FullAdder_29_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_28 = FullAdder_28_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_lo_hi_lo_lo = {mycout_30,mycout_29,mycout_28,mycout_27,mycout_26,mycout_25}; // @[Adder.scala 35:21]
  wire  mycout_33 = FullAdder_33_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_32 = FullAdder_32_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_31 = FullAdder_31_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_36 = FullAdder_36_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_35 = FullAdder_35_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_34 = FullAdder_34_io_cout; // @[Adder.scala 22:20 31:15]
  wire [11:0] io_Cout_lo_hi_lo = {mycout_36,mycout_35,mycout_34,mycout_33,mycout_32,mycout_31,io_Cout_lo_hi_lo_lo}; // @[Adder.scala 35:21]
  wire  mycout_39 = FullAdder_39_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_38 = FullAdder_38_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_37 = FullAdder_37_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_42 = FullAdder_42_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_41 = FullAdder_41_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_40 = FullAdder_40_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_lo_hi_hi_lo = {mycout_42,mycout_41,mycout_40,mycout_39,mycout_38,mycout_37}; // @[Adder.scala 35:21]
  wire  mycout_45 = FullAdder_45_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_44 = FullAdder_44_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_43 = FullAdder_43_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_47 = FullAdder_47_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_46 = FullAdder_46_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_49 = FullAdder_49_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_48 = FullAdder_48_io_cout; // @[Adder.scala 22:20 31:15]
  wire [49:0] io_Cout_lo = {mycout_49,mycout_48,mycout_47,mycout_46,mycout_45,mycout_44,mycout_43,io_Cout_lo_hi_hi_lo,
    io_Cout_lo_hi_lo,io_Cout_lo_lo}; // @[Adder.scala 35:21]
  wire  mycout_52 = FullAdder_52_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_51 = FullAdder_51_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_50 = FullAdder_50_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_55 = FullAdder_55_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_54 = FullAdder_54_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_53 = FullAdder_53_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_hi_lo_lo_lo = {mycout_55,mycout_54,mycout_53,mycout_52,mycout_51,mycout_50}; // @[Adder.scala 35:21]
  wire  mycout_58 = FullAdder_58_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_57 = FullAdder_57_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_56 = FullAdder_56_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_61 = FullAdder_61_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_60 = FullAdder_60_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_59 = FullAdder_59_io_cout; // @[Adder.scala 22:20 31:15]
  wire [11:0] io_Cout_hi_lo_lo = {mycout_61,mycout_60,mycout_59,mycout_58,mycout_57,mycout_56,io_Cout_hi_lo_lo_lo}; // @[Adder.scala 35:21]
  wire  mycout_64 = FullAdder_64_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_63 = FullAdder_63_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_62 = FullAdder_62_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_67 = FullAdder_67_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_66 = FullAdder_66_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_65 = FullAdder_65_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_hi_lo_hi_lo = {mycout_67,mycout_66,mycout_65,mycout_64,mycout_63,mycout_62}; // @[Adder.scala 35:21]
  wire  mycout_70 = FullAdder_70_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_69 = FullAdder_69_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_68 = FullAdder_68_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_72 = FullAdder_72_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_71 = FullAdder_71_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_74 = FullAdder_74_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_73 = FullAdder_73_io_cout; // @[Adder.scala 22:20 31:15]
  wire [24:0] io_Cout_hi_lo = {mycout_74,mycout_73,mycout_72,mycout_71,mycout_70,mycout_69,mycout_68,io_Cout_hi_lo_hi_lo
    ,io_Cout_hi_lo_lo}; // @[Adder.scala 35:21]
  wire  mycout_77 = FullAdder_77_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_76 = FullAdder_76_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_75 = FullAdder_75_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_80 = FullAdder_80_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_79 = FullAdder_79_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_78 = FullAdder_78_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_hi_hi_lo_lo = {mycout_80,mycout_79,mycout_78,mycout_77,mycout_76,mycout_75}; // @[Adder.scala 35:21]
  wire  mycout_83 = FullAdder_83_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_82 = FullAdder_82_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_81 = FullAdder_81_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_86 = FullAdder_86_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_85 = FullAdder_85_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_84 = FullAdder_84_io_cout; // @[Adder.scala 22:20 31:15]
  wire [11:0] io_Cout_hi_hi_lo = {mycout_86,mycout_85,mycout_84,mycout_83,mycout_82,mycout_81,io_Cout_hi_hi_lo_lo}; // @[Adder.scala 35:21]
  wire  mycout_89 = FullAdder_89_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_88 = FullAdder_88_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_87 = FullAdder_87_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_92 = FullAdder_92_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_91 = FullAdder_91_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_90 = FullAdder_90_io_cout; // @[Adder.scala 22:20 31:15]
  wire [5:0] io_Cout_hi_hi_hi_lo = {mycout_92,mycout_91,mycout_90,mycout_89,mycout_88,mycout_87}; // @[Adder.scala 35:21]
  wire  mycout_95 = FullAdder_95_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_94 = FullAdder_94_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_93 = FullAdder_93_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_97 = FullAdder_97_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_96 = FullAdder_96_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_99 = FullAdder_99_io_cout; // @[Adder.scala 22:20 31:15]
  wire  mycout_98 = FullAdder_98_io_cout; // @[Adder.scala 22:20 31:15]
  wire [49:0] io_Cout_hi = {mycout_99,mycout_98,mycout_97,mycout_96,mycout_95,mycout_94,mycout_93,io_Cout_hi_hi_hi_lo,
    io_Cout_hi_hi_lo,io_Cout_hi_lo}; // @[Adder.scala 35:21]
  FullAdder FullAdder ( // @[Adder.scala 19:35]
    .io_a(FullAdder_io_a),
    .io_b(FullAdder_io_b),
    .io_cin(FullAdder_io_cin),
    .io_sum(FullAdder_io_sum),
    .io_cout(FullAdder_io_cout)
  );
  FullAdder FullAdder_1 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_1_io_a),
    .io_b(FullAdder_1_io_b),
    .io_cin(FullAdder_1_io_cin),
    .io_sum(FullAdder_1_io_sum),
    .io_cout(FullAdder_1_io_cout)
  );
  FullAdder FullAdder_2 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_2_io_a),
    .io_b(FullAdder_2_io_b),
    .io_cin(FullAdder_2_io_cin),
    .io_sum(FullAdder_2_io_sum),
    .io_cout(FullAdder_2_io_cout)
  );
  FullAdder FullAdder_3 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_3_io_a),
    .io_b(FullAdder_3_io_b),
    .io_cin(FullAdder_3_io_cin),
    .io_sum(FullAdder_3_io_sum),
    .io_cout(FullAdder_3_io_cout)
  );
  FullAdder FullAdder_4 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_4_io_a),
    .io_b(FullAdder_4_io_b),
    .io_cin(FullAdder_4_io_cin),
    .io_sum(FullAdder_4_io_sum),
    .io_cout(FullAdder_4_io_cout)
  );
  FullAdder FullAdder_5 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_5_io_a),
    .io_b(FullAdder_5_io_b),
    .io_cin(FullAdder_5_io_cin),
    .io_sum(FullAdder_5_io_sum),
    .io_cout(FullAdder_5_io_cout)
  );
  FullAdder FullAdder_6 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_6_io_a),
    .io_b(FullAdder_6_io_b),
    .io_cin(FullAdder_6_io_cin),
    .io_sum(FullAdder_6_io_sum),
    .io_cout(FullAdder_6_io_cout)
  );
  FullAdder FullAdder_7 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_7_io_a),
    .io_b(FullAdder_7_io_b),
    .io_cin(FullAdder_7_io_cin),
    .io_sum(FullAdder_7_io_sum),
    .io_cout(FullAdder_7_io_cout)
  );
  FullAdder FullAdder_8 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_8_io_a),
    .io_b(FullAdder_8_io_b),
    .io_cin(FullAdder_8_io_cin),
    .io_sum(FullAdder_8_io_sum),
    .io_cout(FullAdder_8_io_cout)
  );
  FullAdder FullAdder_9 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_9_io_a),
    .io_b(FullAdder_9_io_b),
    .io_cin(FullAdder_9_io_cin),
    .io_sum(FullAdder_9_io_sum),
    .io_cout(FullAdder_9_io_cout)
  );
  FullAdder FullAdder_10 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_10_io_a),
    .io_b(FullAdder_10_io_b),
    .io_cin(FullAdder_10_io_cin),
    .io_sum(FullAdder_10_io_sum),
    .io_cout(FullAdder_10_io_cout)
  );
  FullAdder FullAdder_11 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_11_io_a),
    .io_b(FullAdder_11_io_b),
    .io_cin(FullAdder_11_io_cin),
    .io_sum(FullAdder_11_io_sum),
    .io_cout(FullAdder_11_io_cout)
  );
  FullAdder FullAdder_12 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_12_io_a),
    .io_b(FullAdder_12_io_b),
    .io_cin(FullAdder_12_io_cin),
    .io_sum(FullAdder_12_io_sum),
    .io_cout(FullAdder_12_io_cout)
  );
  FullAdder FullAdder_13 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_13_io_a),
    .io_b(FullAdder_13_io_b),
    .io_cin(FullAdder_13_io_cin),
    .io_sum(FullAdder_13_io_sum),
    .io_cout(FullAdder_13_io_cout)
  );
  FullAdder FullAdder_14 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_14_io_a),
    .io_b(FullAdder_14_io_b),
    .io_cin(FullAdder_14_io_cin),
    .io_sum(FullAdder_14_io_sum),
    .io_cout(FullAdder_14_io_cout)
  );
  FullAdder FullAdder_15 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_15_io_a),
    .io_b(FullAdder_15_io_b),
    .io_cin(FullAdder_15_io_cin),
    .io_sum(FullAdder_15_io_sum),
    .io_cout(FullAdder_15_io_cout)
  );
  FullAdder FullAdder_16 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_16_io_a),
    .io_b(FullAdder_16_io_b),
    .io_cin(FullAdder_16_io_cin),
    .io_sum(FullAdder_16_io_sum),
    .io_cout(FullAdder_16_io_cout)
  );
  FullAdder FullAdder_17 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_17_io_a),
    .io_b(FullAdder_17_io_b),
    .io_cin(FullAdder_17_io_cin),
    .io_sum(FullAdder_17_io_sum),
    .io_cout(FullAdder_17_io_cout)
  );
  FullAdder FullAdder_18 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_18_io_a),
    .io_b(FullAdder_18_io_b),
    .io_cin(FullAdder_18_io_cin),
    .io_sum(FullAdder_18_io_sum),
    .io_cout(FullAdder_18_io_cout)
  );
  FullAdder FullAdder_19 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_19_io_a),
    .io_b(FullAdder_19_io_b),
    .io_cin(FullAdder_19_io_cin),
    .io_sum(FullAdder_19_io_sum),
    .io_cout(FullAdder_19_io_cout)
  );
  FullAdder FullAdder_20 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_20_io_a),
    .io_b(FullAdder_20_io_b),
    .io_cin(FullAdder_20_io_cin),
    .io_sum(FullAdder_20_io_sum),
    .io_cout(FullAdder_20_io_cout)
  );
  FullAdder FullAdder_21 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_21_io_a),
    .io_b(FullAdder_21_io_b),
    .io_cin(FullAdder_21_io_cin),
    .io_sum(FullAdder_21_io_sum),
    .io_cout(FullAdder_21_io_cout)
  );
  FullAdder FullAdder_22 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_22_io_a),
    .io_b(FullAdder_22_io_b),
    .io_cin(FullAdder_22_io_cin),
    .io_sum(FullAdder_22_io_sum),
    .io_cout(FullAdder_22_io_cout)
  );
  FullAdder FullAdder_23 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_23_io_a),
    .io_b(FullAdder_23_io_b),
    .io_cin(FullAdder_23_io_cin),
    .io_sum(FullAdder_23_io_sum),
    .io_cout(FullAdder_23_io_cout)
  );
  FullAdder FullAdder_24 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_24_io_a),
    .io_b(FullAdder_24_io_b),
    .io_cin(FullAdder_24_io_cin),
    .io_sum(FullAdder_24_io_sum),
    .io_cout(FullAdder_24_io_cout)
  );
  FullAdder FullAdder_25 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_25_io_a),
    .io_b(FullAdder_25_io_b),
    .io_cin(FullAdder_25_io_cin),
    .io_sum(FullAdder_25_io_sum),
    .io_cout(FullAdder_25_io_cout)
  );
  FullAdder FullAdder_26 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_26_io_a),
    .io_b(FullAdder_26_io_b),
    .io_cin(FullAdder_26_io_cin),
    .io_sum(FullAdder_26_io_sum),
    .io_cout(FullAdder_26_io_cout)
  );
  FullAdder FullAdder_27 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_27_io_a),
    .io_b(FullAdder_27_io_b),
    .io_cin(FullAdder_27_io_cin),
    .io_sum(FullAdder_27_io_sum),
    .io_cout(FullAdder_27_io_cout)
  );
  FullAdder FullAdder_28 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_28_io_a),
    .io_b(FullAdder_28_io_b),
    .io_cin(FullAdder_28_io_cin),
    .io_sum(FullAdder_28_io_sum),
    .io_cout(FullAdder_28_io_cout)
  );
  FullAdder FullAdder_29 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_29_io_a),
    .io_b(FullAdder_29_io_b),
    .io_cin(FullAdder_29_io_cin),
    .io_sum(FullAdder_29_io_sum),
    .io_cout(FullAdder_29_io_cout)
  );
  FullAdder FullAdder_30 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_30_io_a),
    .io_b(FullAdder_30_io_b),
    .io_cin(FullAdder_30_io_cin),
    .io_sum(FullAdder_30_io_sum),
    .io_cout(FullAdder_30_io_cout)
  );
  FullAdder FullAdder_31 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_31_io_a),
    .io_b(FullAdder_31_io_b),
    .io_cin(FullAdder_31_io_cin),
    .io_sum(FullAdder_31_io_sum),
    .io_cout(FullAdder_31_io_cout)
  );
  FullAdder FullAdder_32 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_32_io_a),
    .io_b(FullAdder_32_io_b),
    .io_cin(FullAdder_32_io_cin),
    .io_sum(FullAdder_32_io_sum),
    .io_cout(FullAdder_32_io_cout)
  );
  FullAdder FullAdder_33 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_33_io_a),
    .io_b(FullAdder_33_io_b),
    .io_cin(FullAdder_33_io_cin),
    .io_sum(FullAdder_33_io_sum),
    .io_cout(FullAdder_33_io_cout)
  );
  FullAdder FullAdder_34 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_34_io_a),
    .io_b(FullAdder_34_io_b),
    .io_cin(FullAdder_34_io_cin),
    .io_sum(FullAdder_34_io_sum),
    .io_cout(FullAdder_34_io_cout)
  );
  FullAdder FullAdder_35 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_35_io_a),
    .io_b(FullAdder_35_io_b),
    .io_cin(FullAdder_35_io_cin),
    .io_sum(FullAdder_35_io_sum),
    .io_cout(FullAdder_35_io_cout)
  );
  FullAdder FullAdder_36 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_36_io_a),
    .io_b(FullAdder_36_io_b),
    .io_cin(FullAdder_36_io_cin),
    .io_sum(FullAdder_36_io_sum),
    .io_cout(FullAdder_36_io_cout)
  );
  FullAdder FullAdder_37 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_37_io_a),
    .io_b(FullAdder_37_io_b),
    .io_cin(FullAdder_37_io_cin),
    .io_sum(FullAdder_37_io_sum),
    .io_cout(FullAdder_37_io_cout)
  );
  FullAdder FullAdder_38 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_38_io_a),
    .io_b(FullAdder_38_io_b),
    .io_cin(FullAdder_38_io_cin),
    .io_sum(FullAdder_38_io_sum),
    .io_cout(FullAdder_38_io_cout)
  );
  FullAdder FullAdder_39 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_39_io_a),
    .io_b(FullAdder_39_io_b),
    .io_cin(FullAdder_39_io_cin),
    .io_sum(FullAdder_39_io_sum),
    .io_cout(FullAdder_39_io_cout)
  );
  FullAdder FullAdder_40 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_40_io_a),
    .io_b(FullAdder_40_io_b),
    .io_cin(FullAdder_40_io_cin),
    .io_sum(FullAdder_40_io_sum),
    .io_cout(FullAdder_40_io_cout)
  );
  FullAdder FullAdder_41 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_41_io_a),
    .io_b(FullAdder_41_io_b),
    .io_cin(FullAdder_41_io_cin),
    .io_sum(FullAdder_41_io_sum),
    .io_cout(FullAdder_41_io_cout)
  );
  FullAdder FullAdder_42 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_42_io_a),
    .io_b(FullAdder_42_io_b),
    .io_cin(FullAdder_42_io_cin),
    .io_sum(FullAdder_42_io_sum),
    .io_cout(FullAdder_42_io_cout)
  );
  FullAdder FullAdder_43 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_43_io_a),
    .io_b(FullAdder_43_io_b),
    .io_cin(FullAdder_43_io_cin),
    .io_sum(FullAdder_43_io_sum),
    .io_cout(FullAdder_43_io_cout)
  );
  FullAdder FullAdder_44 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_44_io_a),
    .io_b(FullAdder_44_io_b),
    .io_cin(FullAdder_44_io_cin),
    .io_sum(FullAdder_44_io_sum),
    .io_cout(FullAdder_44_io_cout)
  );
  FullAdder FullAdder_45 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_45_io_a),
    .io_b(FullAdder_45_io_b),
    .io_cin(FullAdder_45_io_cin),
    .io_sum(FullAdder_45_io_sum),
    .io_cout(FullAdder_45_io_cout)
  );
  FullAdder FullAdder_46 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_46_io_a),
    .io_b(FullAdder_46_io_b),
    .io_cin(FullAdder_46_io_cin),
    .io_sum(FullAdder_46_io_sum),
    .io_cout(FullAdder_46_io_cout)
  );
  FullAdder FullAdder_47 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_47_io_a),
    .io_b(FullAdder_47_io_b),
    .io_cin(FullAdder_47_io_cin),
    .io_sum(FullAdder_47_io_sum),
    .io_cout(FullAdder_47_io_cout)
  );
  FullAdder FullAdder_48 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_48_io_a),
    .io_b(FullAdder_48_io_b),
    .io_cin(FullAdder_48_io_cin),
    .io_sum(FullAdder_48_io_sum),
    .io_cout(FullAdder_48_io_cout)
  );
  FullAdder FullAdder_49 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_49_io_a),
    .io_b(FullAdder_49_io_b),
    .io_cin(FullAdder_49_io_cin),
    .io_sum(FullAdder_49_io_sum),
    .io_cout(FullAdder_49_io_cout)
  );
  FullAdder FullAdder_50 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_50_io_a),
    .io_b(FullAdder_50_io_b),
    .io_cin(FullAdder_50_io_cin),
    .io_sum(FullAdder_50_io_sum),
    .io_cout(FullAdder_50_io_cout)
  );
  FullAdder FullAdder_51 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_51_io_a),
    .io_b(FullAdder_51_io_b),
    .io_cin(FullAdder_51_io_cin),
    .io_sum(FullAdder_51_io_sum),
    .io_cout(FullAdder_51_io_cout)
  );
  FullAdder FullAdder_52 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_52_io_a),
    .io_b(FullAdder_52_io_b),
    .io_cin(FullAdder_52_io_cin),
    .io_sum(FullAdder_52_io_sum),
    .io_cout(FullAdder_52_io_cout)
  );
  FullAdder FullAdder_53 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_53_io_a),
    .io_b(FullAdder_53_io_b),
    .io_cin(FullAdder_53_io_cin),
    .io_sum(FullAdder_53_io_sum),
    .io_cout(FullAdder_53_io_cout)
  );
  FullAdder FullAdder_54 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_54_io_a),
    .io_b(FullAdder_54_io_b),
    .io_cin(FullAdder_54_io_cin),
    .io_sum(FullAdder_54_io_sum),
    .io_cout(FullAdder_54_io_cout)
  );
  FullAdder FullAdder_55 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_55_io_a),
    .io_b(FullAdder_55_io_b),
    .io_cin(FullAdder_55_io_cin),
    .io_sum(FullAdder_55_io_sum),
    .io_cout(FullAdder_55_io_cout)
  );
  FullAdder FullAdder_56 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_56_io_a),
    .io_b(FullAdder_56_io_b),
    .io_cin(FullAdder_56_io_cin),
    .io_sum(FullAdder_56_io_sum),
    .io_cout(FullAdder_56_io_cout)
  );
  FullAdder FullAdder_57 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_57_io_a),
    .io_b(FullAdder_57_io_b),
    .io_cin(FullAdder_57_io_cin),
    .io_sum(FullAdder_57_io_sum),
    .io_cout(FullAdder_57_io_cout)
  );
  FullAdder FullAdder_58 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_58_io_a),
    .io_b(FullAdder_58_io_b),
    .io_cin(FullAdder_58_io_cin),
    .io_sum(FullAdder_58_io_sum),
    .io_cout(FullAdder_58_io_cout)
  );
  FullAdder FullAdder_59 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_59_io_a),
    .io_b(FullAdder_59_io_b),
    .io_cin(FullAdder_59_io_cin),
    .io_sum(FullAdder_59_io_sum),
    .io_cout(FullAdder_59_io_cout)
  );
  FullAdder FullAdder_60 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_60_io_a),
    .io_b(FullAdder_60_io_b),
    .io_cin(FullAdder_60_io_cin),
    .io_sum(FullAdder_60_io_sum),
    .io_cout(FullAdder_60_io_cout)
  );
  FullAdder FullAdder_61 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_61_io_a),
    .io_b(FullAdder_61_io_b),
    .io_cin(FullAdder_61_io_cin),
    .io_sum(FullAdder_61_io_sum),
    .io_cout(FullAdder_61_io_cout)
  );
  FullAdder FullAdder_62 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_62_io_a),
    .io_b(FullAdder_62_io_b),
    .io_cin(FullAdder_62_io_cin),
    .io_sum(FullAdder_62_io_sum),
    .io_cout(FullAdder_62_io_cout)
  );
  FullAdder FullAdder_63 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_63_io_a),
    .io_b(FullAdder_63_io_b),
    .io_cin(FullAdder_63_io_cin),
    .io_sum(FullAdder_63_io_sum),
    .io_cout(FullAdder_63_io_cout)
  );
  FullAdder FullAdder_64 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_64_io_a),
    .io_b(FullAdder_64_io_b),
    .io_cin(FullAdder_64_io_cin),
    .io_sum(FullAdder_64_io_sum),
    .io_cout(FullAdder_64_io_cout)
  );
  FullAdder FullAdder_65 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_65_io_a),
    .io_b(FullAdder_65_io_b),
    .io_cin(FullAdder_65_io_cin),
    .io_sum(FullAdder_65_io_sum),
    .io_cout(FullAdder_65_io_cout)
  );
  FullAdder FullAdder_66 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_66_io_a),
    .io_b(FullAdder_66_io_b),
    .io_cin(FullAdder_66_io_cin),
    .io_sum(FullAdder_66_io_sum),
    .io_cout(FullAdder_66_io_cout)
  );
  FullAdder FullAdder_67 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_67_io_a),
    .io_b(FullAdder_67_io_b),
    .io_cin(FullAdder_67_io_cin),
    .io_sum(FullAdder_67_io_sum),
    .io_cout(FullAdder_67_io_cout)
  );
  FullAdder FullAdder_68 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_68_io_a),
    .io_b(FullAdder_68_io_b),
    .io_cin(FullAdder_68_io_cin),
    .io_sum(FullAdder_68_io_sum),
    .io_cout(FullAdder_68_io_cout)
  );
  FullAdder FullAdder_69 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_69_io_a),
    .io_b(FullAdder_69_io_b),
    .io_cin(FullAdder_69_io_cin),
    .io_sum(FullAdder_69_io_sum),
    .io_cout(FullAdder_69_io_cout)
  );
  FullAdder FullAdder_70 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_70_io_a),
    .io_b(FullAdder_70_io_b),
    .io_cin(FullAdder_70_io_cin),
    .io_sum(FullAdder_70_io_sum),
    .io_cout(FullAdder_70_io_cout)
  );
  FullAdder FullAdder_71 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_71_io_a),
    .io_b(FullAdder_71_io_b),
    .io_cin(FullAdder_71_io_cin),
    .io_sum(FullAdder_71_io_sum),
    .io_cout(FullAdder_71_io_cout)
  );
  FullAdder FullAdder_72 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_72_io_a),
    .io_b(FullAdder_72_io_b),
    .io_cin(FullAdder_72_io_cin),
    .io_sum(FullAdder_72_io_sum),
    .io_cout(FullAdder_72_io_cout)
  );
  FullAdder FullAdder_73 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_73_io_a),
    .io_b(FullAdder_73_io_b),
    .io_cin(FullAdder_73_io_cin),
    .io_sum(FullAdder_73_io_sum),
    .io_cout(FullAdder_73_io_cout)
  );
  FullAdder FullAdder_74 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_74_io_a),
    .io_b(FullAdder_74_io_b),
    .io_cin(FullAdder_74_io_cin),
    .io_sum(FullAdder_74_io_sum),
    .io_cout(FullAdder_74_io_cout)
  );
  FullAdder FullAdder_75 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_75_io_a),
    .io_b(FullAdder_75_io_b),
    .io_cin(FullAdder_75_io_cin),
    .io_sum(FullAdder_75_io_sum),
    .io_cout(FullAdder_75_io_cout)
  );
  FullAdder FullAdder_76 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_76_io_a),
    .io_b(FullAdder_76_io_b),
    .io_cin(FullAdder_76_io_cin),
    .io_sum(FullAdder_76_io_sum),
    .io_cout(FullAdder_76_io_cout)
  );
  FullAdder FullAdder_77 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_77_io_a),
    .io_b(FullAdder_77_io_b),
    .io_cin(FullAdder_77_io_cin),
    .io_sum(FullAdder_77_io_sum),
    .io_cout(FullAdder_77_io_cout)
  );
  FullAdder FullAdder_78 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_78_io_a),
    .io_b(FullAdder_78_io_b),
    .io_cin(FullAdder_78_io_cin),
    .io_sum(FullAdder_78_io_sum),
    .io_cout(FullAdder_78_io_cout)
  );
  FullAdder FullAdder_79 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_79_io_a),
    .io_b(FullAdder_79_io_b),
    .io_cin(FullAdder_79_io_cin),
    .io_sum(FullAdder_79_io_sum),
    .io_cout(FullAdder_79_io_cout)
  );
  FullAdder FullAdder_80 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_80_io_a),
    .io_b(FullAdder_80_io_b),
    .io_cin(FullAdder_80_io_cin),
    .io_sum(FullAdder_80_io_sum),
    .io_cout(FullAdder_80_io_cout)
  );
  FullAdder FullAdder_81 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_81_io_a),
    .io_b(FullAdder_81_io_b),
    .io_cin(FullAdder_81_io_cin),
    .io_sum(FullAdder_81_io_sum),
    .io_cout(FullAdder_81_io_cout)
  );
  FullAdder FullAdder_82 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_82_io_a),
    .io_b(FullAdder_82_io_b),
    .io_cin(FullAdder_82_io_cin),
    .io_sum(FullAdder_82_io_sum),
    .io_cout(FullAdder_82_io_cout)
  );
  FullAdder FullAdder_83 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_83_io_a),
    .io_b(FullAdder_83_io_b),
    .io_cin(FullAdder_83_io_cin),
    .io_sum(FullAdder_83_io_sum),
    .io_cout(FullAdder_83_io_cout)
  );
  FullAdder FullAdder_84 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_84_io_a),
    .io_b(FullAdder_84_io_b),
    .io_cin(FullAdder_84_io_cin),
    .io_sum(FullAdder_84_io_sum),
    .io_cout(FullAdder_84_io_cout)
  );
  FullAdder FullAdder_85 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_85_io_a),
    .io_b(FullAdder_85_io_b),
    .io_cin(FullAdder_85_io_cin),
    .io_sum(FullAdder_85_io_sum),
    .io_cout(FullAdder_85_io_cout)
  );
  FullAdder FullAdder_86 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_86_io_a),
    .io_b(FullAdder_86_io_b),
    .io_cin(FullAdder_86_io_cin),
    .io_sum(FullAdder_86_io_sum),
    .io_cout(FullAdder_86_io_cout)
  );
  FullAdder FullAdder_87 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_87_io_a),
    .io_b(FullAdder_87_io_b),
    .io_cin(FullAdder_87_io_cin),
    .io_sum(FullAdder_87_io_sum),
    .io_cout(FullAdder_87_io_cout)
  );
  FullAdder FullAdder_88 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_88_io_a),
    .io_b(FullAdder_88_io_b),
    .io_cin(FullAdder_88_io_cin),
    .io_sum(FullAdder_88_io_sum),
    .io_cout(FullAdder_88_io_cout)
  );
  FullAdder FullAdder_89 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_89_io_a),
    .io_b(FullAdder_89_io_b),
    .io_cin(FullAdder_89_io_cin),
    .io_sum(FullAdder_89_io_sum),
    .io_cout(FullAdder_89_io_cout)
  );
  FullAdder FullAdder_90 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_90_io_a),
    .io_b(FullAdder_90_io_b),
    .io_cin(FullAdder_90_io_cin),
    .io_sum(FullAdder_90_io_sum),
    .io_cout(FullAdder_90_io_cout)
  );
  FullAdder FullAdder_91 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_91_io_a),
    .io_b(FullAdder_91_io_b),
    .io_cin(FullAdder_91_io_cin),
    .io_sum(FullAdder_91_io_sum),
    .io_cout(FullAdder_91_io_cout)
  );
  FullAdder FullAdder_92 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_92_io_a),
    .io_b(FullAdder_92_io_b),
    .io_cin(FullAdder_92_io_cin),
    .io_sum(FullAdder_92_io_sum),
    .io_cout(FullAdder_92_io_cout)
  );
  FullAdder FullAdder_93 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_93_io_a),
    .io_b(FullAdder_93_io_b),
    .io_cin(FullAdder_93_io_cin),
    .io_sum(FullAdder_93_io_sum),
    .io_cout(FullAdder_93_io_cout)
  );
  FullAdder FullAdder_94 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_94_io_a),
    .io_b(FullAdder_94_io_b),
    .io_cin(FullAdder_94_io_cin),
    .io_sum(FullAdder_94_io_sum),
    .io_cout(FullAdder_94_io_cout)
  );
  FullAdder FullAdder_95 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_95_io_a),
    .io_b(FullAdder_95_io_b),
    .io_cin(FullAdder_95_io_cin),
    .io_sum(FullAdder_95_io_sum),
    .io_cout(FullAdder_95_io_cout)
  );
  FullAdder FullAdder_96 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_96_io_a),
    .io_b(FullAdder_96_io_b),
    .io_cin(FullAdder_96_io_cin),
    .io_sum(FullAdder_96_io_sum),
    .io_cout(FullAdder_96_io_cout)
  );
  FullAdder FullAdder_97 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_97_io_a),
    .io_b(FullAdder_97_io_b),
    .io_cin(FullAdder_97_io_cin),
    .io_sum(FullAdder_97_io_sum),
    .io_cout(FullAdder_97_io_cout)
  );
  FullAdder FullAdder_98 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_98_io_a),
    .io_b(FullAdder_98_io_b),
    .io_cin(FullAdder_98_io_cin),
    .io_sum(FullAdder_98_io_sum),
    .io_cout(FullAdder_98_io_cout)
  );
  FullAdder FullAdder_99 ( // @[Adder.scala 19:35]
    .io_a(FullAdder_99_io_a),
    .io_b(FullAdder_99_io_b),
    .io_cin(FullAdder_99_io_cin),
    .io_sum(FullAdder_99_io_sum),
    .io_cout(FullAdder_99_io_cout)
  );
  assign io_Sum = {io_Sum_hi,io_Sum_lo}; // @[Adder.scala 34:17]
  assign io_Cout = {io_Cout_hi,io_Cout_lo}; // @[Adder.scala 35:21]
  assign FullAdder_io_a = io_A[0]; // @[Adder.scala 27:21]
  assign FullAdder_io_b = io_B[0]; // @[Adder.scala 28:21]
  assign FullAdder_io_cin = io_Cin; // @[Adder.scala 20:19 24:12]
  assign FullAdder_1_io_a = io_A[1]; // @[Adder.scala 27:21]
  assign FullAdder_1_io_b = io_B[1]; // @[Adder.scala 28:21]
  assign FullAdder_1_io_cin = FullAdder_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_2_io_a = io_A[2]; // @[Adder.scala 27:21]
  assign FullAdder_2_io_b = io_B[2]; // @[Adder.scala 28:21]
  assign FullAdder_2_io_cin = FullAdder_1_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_3_io_a = io_A[3]; // @[Adder.scala 27:21]
  assign FullAdder_3_io_b = io_B[3]; // @[Adder.scala 28:21]
  assign FullAdder_3_io_cin = FullAdder_2_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_4_io_a = io_A[4]; // @[Adder.scala 27:21]
  assign FullAdder_4_io_b = io_B[4]; // @[Adder.scala 28:21]
  assign FullAdder_4_io_cin = FullAdder_3_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_5_io_a = io_A[5]; // @[Adder.scala 27:21]
  assign FullAdder_5_io_b = io_B[5]; // @[Adder.scala 28:21]
  assign FullAdder_5_io_cin = FullAdder_4_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_6_io_a = io_A[6]; // @[Adder.scala 27:21]
  assign FullAdder_6_io_b = io_B[6]; // @[Adder.scala 28:21]
  assign FullAdder_6_io_cin = FullAdder_5_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_7_io_a = io_A[7]; // @[Adder.scala 27:21]
  assign FullAdder_7_io_b = io_B[7]; // @[Adder.scala 28:21]
  assign FullAdder_7_io_cin = FullAdder_6_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_8_io_a = io_A[8]; // @[Adder.scala 27:21]
  assign FullAdder_8_io_b = io_B[8]; // @[Adder.scala 28:21]
  assign FullAdder_8_io_cin = FullAdder_7_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_9_io_a = io_A[9]; // @[Adder.scala 27:21]
  assign FullAdder_9_io_b = io_B[9]; // @[Adder.scala 28:21]
  assign FullAdder_9_io_cin = FullAdder_8_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_10_io_a = io_A[10]; // @[Adder.scala 27:21]
  assign FullAdder_10_io_b = io_B[10]; // @[Adder.scala 28:21]
  assign FullAdder_10_io_cin = FullAdder_9_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_11_io_a = io_A[11]; // @[Adder.scala 27:21]
  assign FullAdder_11_io_b = io_B[11]; // @[Adder.scala 28:21]
  assign FullAdder_11_io_cin = FullAdder_10_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_12_io_a = io_A[12]; // @[Adder.scala 27:21]
  assign FullAdder_12_io_b = io_B[12]; // @[Adder.scala 28:21]
  assign FullAdder_12_io_cin = FullAdder_11_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_13_io_a = io_A[13]; // @[Adder.scala 27:21]
  assign FullAdder_13_io_b = io_B[13]; // @[Adder.scala 28:21]
  assign FullAdder_13_io_cin = FullAdder_12_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_14_io_a = io_A[14]; // @[Adder.scala 27:21]
  assign FullAdder_14_io_b = io_B[14]; // @[Adder.scala 28:21]
  assign FullAdder_14_io_cin = FullAdder_13_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_15_io_a = io_A[15]; // @[Adder.scala 27:21]
  assign FullAdder_15_io_b = io_B[15]; // @[Adder.scala 28:21]
  assign FullAdder_15_io_cin = FullAdder_14_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_16_io_a = io_A[16]; // @[Adder.scala 27:21]
  assign FullAdder_16_io_b = io_B[16]; // @[Adder.scala 28:21]
  assign FullAdder_16_io_cin = FullAdder_15_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_17_io_a = io_A[17]; // @[Adder.scala 27:21]
  assign FullAdder_17_io_b = io_B[17]; // @[Adder.scala 28:21]
  assign FullAdder_17_io_cin = FullAdder_16_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_18_io_a = io_A[18]; // @[Adder.scala 27:21]
  assign FullAdder_18_io_b = io_B[18]; // @[Adder.scala 28:21]
  assign FullAdder_18_io_cin = FullAdder_17_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_19_io_a = io_A[19]; // @[Adder.scala 27:21]
  assign FullAdder_19_io_b = io_B[19]; // @[Adder.scala 28:21]
  assign FullAdder_19_io_cin = FullAdder_18_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_20_io_a = io_A[20]; // @[Adder.scala 27:21]
  assign FullAdder_20_io_b = io_B[20]; // @[Adder.scala 28:21]
  assign FullAdder_20_io_cin = FullAdder_19_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_21_io_a = io_A[21]; // @[Adder.scala 27:21]
  assign FullAdder_21_io_b = io_B[21]; // @[Adder.scala 28:21]
  assign FullAdder_21_io_cin = FullAdder_20_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_22_io_a = io_A[22]; // @[Adder.scala 27:21]
  assign FullAdder_22_io_b = io_B[22]; // @[Adder.scala 28:21]
  assign FullAdder_22_io_cin = FullAdder_21_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_23_io_a = io_A[23]; // @[Adder.scala 27:21]
  assign FullAdder_23_io_b = io_B[23]; // @[Adder.scala 28:21]
  assign FullAdder_23_io_cin = FullAdder_22_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_24_io_a = io_A[24]; // @[Adder.scala 27:21]
  assign FullAdder_24_io_b = io_B[24]; // @[Adder.scala 28:21]
  assign FullAdder_24_io_cin = FullAdder_23_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_25_io_a = io_A[25]; // @[Adder.scala 27:21]
  assign FullAdder_25_io_b = io_B[25]; // @[Adder.scala 28:21]
  assign FullAdder_25_io_cin = FullAdder_24_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_26_io_a = io_A[26]; // @[Adder.scala 27:21]
  assign FullAdder_26_io_b = io_B[26]; // @[Adder.scala 28:21]
  assign FullAdder_26_io_cin = FullAdder_25_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_27_io_a = io_A[27]; // @[Adder.scala 27:21]
  assign FullAdder_27_io_b = io_B[27]; // @[Adder.scala 28:21]
  assign FullAdder_27_io_cin = FullAdder_26_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_28_io_a = io_A[28]; // @[Adder.scala 27:21]
  assign FullAdder_28_io_b = io_B[28]; // @[Adder.scala 28:21]
  assign FullAdder_28_io_cin = FullAdder_27_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_29_io_a = io_A[29]; // @[Adder.scala 27:21]
  assign FullAdder_29_io_b = io_B[29]; // @[Adder.scala 28:21]
  assign FullAdder_29_io_cin = FullAdder_28_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_30_io_a = io_A[30]; // @[Adder.scala 27:21]
  assign FullAdder_30_io_b = io_B[30]; // @[Adder.scala 28:21]
  assign FullAdder_30_io_cin = FullAdder_29_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_31_io_a = io_A[31]; // @[Adder.scala 27:21]
  assign FullAdder_31_io_b = io_B[31]; // @[Adder.scala 28:21]
  assign FullAdder_31_io_cin = FullAdder_30_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_32_io_a = io_A[32]; // @[Adder.scala 27:21]
  assign FullAdder_32_io_b = io_B[32]; // @[Adder.scala 28:21]
  assign FullAdder_32_io_cin = FullAdder_31_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_33_io_a = io_A[33]; // @[Adder.scala 27:21]
  assign FullAdder_33_io_b = io_B[33]; // @[Adder.scala 28:21]
  assign FullAdder_33_io_cin = FullAdder_32_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_34_io_a = io_A[34]; // @[Adder.scala 27:21]
  assign FullAdder_34_io_b = io_B[34]; // @[Adder.scala 28:21]
  assign FullAdder_34_io_cin = FullAdder_33_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_35_io_a = io_A[35]; // @[Adder.scala 27:21]
  assign FullAdder_35_io_b = io_B[35]; // @[Adder.scala 28:21]
  assign FullAdder_35_io_cin = FullAdder_34_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_36_io_a = io_A[36]; // @[Adder.scala 27:21]
  assign FullAdder_36_io_b = io_B[36]; // @[Adder.scala 28:21]
  assign FullAdder_36_io_cin = FullAdder_35_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_37_io_a = io_A[37]; // @[Adder.scala 27:21]
  assign FullAdder_37_io_b = io_B[37]; // @[Adder.scala 28:21]
  assign FullAdder_37_io_cin = FullAdder_36_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_38_io_a = io_A[38]; // @[Adder.scala 27:21]
  assign FullAdder_38_io_b = io_B[38]; // @[Adder.scala 28:21]
  assign FullAdder_38_io_cin = FullAdder_37_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_39_io_a = io_A[39]; // @[Adder.scala 27:21]
  assign FullAdder_39_io_b = io_B[39]; // @[Adder.scala 28:21]
  assign FullAdder_39_io_cin = FullAdder_38_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_40_io_a = io_A[40]; // @[Adder.scala 27:21]
  assign FullAdder_40_io_b = io_B[40]; // @[Adder.scala 28:21]
  assign FullAdder_40_io_cin = FullAdder_39_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_41_io_a = io_A[41]; // @[Adder.scala 27:21]
  assign FullAdder_41_io_b = io_B[41]; // @[Adder.scala 28:21]
  assign FullAdder_41_io_cin = FullAdder_40_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_42_io_a = io_A[42]; // @[Adder.scala 27:21]
  assign FullAdder_42_io_b = io_B[42]; // @[Adder.scala 28:21]
  assign FullAdder_42_io_cin = FullAdder_41_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_43_io_a = io_A[43]; // @[Adder.scala 27:21]
  assign FullAdder_43_io_b = io_B[43]; // @[Adder.scala 28:21]
  assign FullAdder_43_io_cin = FullAdder_42_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_44_io_a = io_A[44]; // @[Adder.scala 27:21]
  assign FullAdder_44_io_b = io_B[44]; // @[Adder.scala 28:21]
  assign FullAdder_44_io_cin = FullAdder_43_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_45_io_a = io_A[45]; // @[Adder.scala 27:21]
  assign FullAdder_45_io_b = io_B[45]; // @[Adder.scala 28:21]
  assign FullAdder_45_io_cin = FullAdder_44_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_46_io_a = io_A[46]; // @[Adder.scala 27:21]
  assign FullAdder_46_io_b = io_B[46]; // @[Adder.scala 28:21]
  assign FullAdder_46_io_cin = FullAdder_45_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_47_io_a = io_A[47]; // @[Adder.scala 27:21]
  assign FullAdder_47_io_b = io_B[47]; // @[Adder.scala 28:21]
  assign FullAdder_47_io_cin = FullAdder_46_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_48_io_a = io_A[48]; // @[Adder.scala 27:21]
  assign FullAdder_48_io_b = io_B[48]; // @[Adder.scala 28:21]
  assign FullAdder_48_io_cin = FullAdder_47_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_49_io_a = io_A[49]; // @[Adder.scala 27:21]
  assign FullAdder_49_io_b = io_B[49]; // @[Adder.scala 28:21]
  assign FullAdder_49_io_cin = FullAdder_48_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_50_io_a = io_A[50]; // @[Adder.scala 27:21]
  assign FullAdder_50_io_b = io_B[50]; // @[Adder.scala 28:21]
  assign FullAdder_50_io_cin = FullAdder_49_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_51_io_a = io_A[51]; // @[Adder.scala 27:21]
  assign FullAdder_51_io_b = io_B[51]; // @[Adder.scala 28:21]
  assign FullAdder_51_io_cin = FullAdder_50_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_52_io_a = io_A[52]; // @[Adder.scala 27:21]
  assign FullAdder_52_io_b = io_B[52]; // @[Adder.scala 28:21]
  assign FullAdder_52_io_cin = FullAdder_51_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_53_io_a = io_A[53]; // @[Adder.scala 27:21]
  assign FullAdder_53_io_b = io_B[53]; // @[Adder.scala 28:21]
  assign FullAdder_53_io_cin = FullAdder_52_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_54_io_a = io_A[54]; // @[Adder.scala 27:21]
  assign FullAdder_54_io_b = io_B[54]; // @[Adder.scala 28:21]
  assign FullAdder_54_io_cin = FullAdder_53_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_55_io_a = io_A[55]; // @[Adder.scala 27:21]
  assign FullAdder_55_io_b = io_B[55]; // @[Adder.scala 28:21]
  assign FullAdder_55_io_cin = FullAdder_54_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_56_io_a = io_A[56]; // @[Adder.scala 27:21]
  assign FullAdder_56_io_b = io_B[56]; // @[Adder.scala 28:21]
  assign FullAdder_56_io_cin = FullAdder_55_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_57_io_a = io_A[57]; // @[Adder.scala 27:21]
  assign FullAdder_57_io_b = io_B[57]; // @[Adder.scala 28:21]
  assign FullAdder_57_io_cin = FullAdder_56_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_58_io_a = io_A[58]; // @[Adder.scala 27:21]
  assign FullAdder_58_io_b = io_B[58]; // @[Adder.scala 28:21]
  assign FullAdder_58_io_cin = FullAdder_57_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_59_io_a = io_A[59]; // @[Adder.scala 27:21]
  assign FullAdder_59_io_b = io_B[59]; // @[Adder.scala 28:21]
  assign FullAdder_59_io_cin = FullAdder_58_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_60_io_a = io_A[60]; // @[Adder.scala 27:21]
  assign FullAdder_60_io_b = io_B[60]; // @[Adder.scala 28:21]
  assign FullAdder_60_io_cin = FullAdder_59_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_61_io_a = io_A[61]; // @[Adder.scala 27:21]
  assign FullAdder_61_io_b = io_B[61]; // @[Adder.scala 28:21]
  assign FullAdder_61_io_cin = FullAdder_60_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_62_io_a = io_A[62]; // @[Adder.scala 27:21]
  assign FullAdder_62_io_b = io_B[62]; // @[Adder.scala 28:21]
  assign FullAdder_62_io_cin = FullAdder_61_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_63_io_a = io_A[63]; // @[Adder.scala 27:21]
  assign FullAdder_63_io_b = io_B[63]; // @[Adder.scala 28:21]
  assign FullAdder_63_io_cin = FullAdder_62_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_64_io_a = io_A[64]; // @[Adder.scala 27:21]
  assign FullAdder_64_io_b = io_B[64]; // @[Adder.scala 28:21]
  assign FullAdder_64_io_cin = FullAdder_63_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_65_io_a = io_A[65]; // @[Adder.scala 27:21]
  assign FullAdder_65_io_b = io_B[65]; // @[Adder.scala 28:21]
  assign FullAdder_65_io_cin = FullAdder_64_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_66_io_a = io_A[66]; // @[Adder.scala 27:21]
  assign FullAdder_66_io_b = io_B[66]; // @[Adder.scala 28:21]
  assign FullAdder_66_io_cin = FullAdder_65_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_67_io_a = io_A[67]; // @[Adder.scala 27:21]
  assign FullAdder_67_io_b = io_B[67]; // @[Adder.scala 28:21]
  assign FullAdder_67_io_cin = FullAdder_66_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_68_io_a = io_A[68]; // @[Adder.scala 27:21]
  assign FullAdder_68_io_b = io_B[68]; // @[Adder.scala 28:21]
  assign FullAdder_68_io_cin = FullAdder_67_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_69_io_a = io_A[69]; // @[Adder.scala 27:21]
  assign FullAdder_69_io_b = io_B[69]; // @[Adder.scala 28:21]
  assign FullAdder_69_io_cin = FullAdder_68_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_70_io_a = io_A[70]; // @[Adder.scala 27:21]
  assign FullAdder_70_io_b = io_B[70]; // @[Adder.scala 28:21]
  assign FullAdder_70_io_cin = FullAdder_69_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_71_io_a = io_A[71]; // @[Adder.scala 27:21]
  assign FullAdder_71_io_b = io_B[71]; // @[Adder.scala 28:21]
  assign FullAdder_71_io_cin = FullAdder_70_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_72_io_a = io_A[72]; // @[Adder.scala 27:21]
  assign FullAdder_72_io_b = io_B[72]; // @[Adder.scala 28:21]
  assign FullAdder_72_io_cin = FullAdder_71_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_73_io_a = io_A[73]; // @[Adder.scala 27:21]
  assign FullAdder_73_io_b = io_B[73]; // @[Adder.scala 28:21]
  assign FullAdder_73_io_cin = FullAdder_72_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_74_io_a = io_A[74]; // @[Adder.scala 27:21]
  assign FullAdder_74_io_b = io_B[74]; // @[Adder.scala 28:21]
  assign FullAdder_74_io_cin = FullAdder_73_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_75_io_a = io_A[75]; // @[Adder.scala 27:21]
  assign FullAdder_75_io_b = io_B[75]; // @[Adder.scala 28:21]
  assign FullAdder_75_io_cin = FullAdder_74_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_76_io_a = io_A[76]; // @[Adder.scala 27:21]
  assign FullAdder_76_io_b = io_B[76]; // @[Adder.scala 28:21]
  assign FullAdder_76_io_cin = FullAdder_75_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_77_io_a = io_A[77]; // @[Adder.scala 27:21]
  assign FullAdder_77_io_b = io_B[77]; // @[Adder.scala 28:21]
  assign FullAdder_77_io_cin = FullAdder_76_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_78_io_a = io_A[78]; // @[Adder.scala 27:21]
  assign FullAdder_78_io_b = io_B[78]; // @[Adder.scala 28:21]
  assign FullAdder_78_io_cin = FullAdder_77_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_79_io_a = io_A[79]; // @[Adder.scala 27:21]
  assign FullAdder_79_io_b = io_B[79]; // @[Adder.scala 28:21]
  assign FullAdder_79_io_cin = FullAdder_78_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_80_io_a = io_A[80]; // @[Adder.scala 27:21]
  assign FullAdder_80_io_b = io_B[80]; // @[Adder.scala 28:21]
  assign FullAdder_80_io_cin = FullAdder_79_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_81_io_a = io_A[81]; // @[Adder.scala 27:21]
  assign FullAdder_81_io_b = io_B[81]; // @[Adder.scala 28:21]
  assign FullAdder_81_io_cin = FullAdder_80_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_82_io_a = io_A[82]; // @[Adder.scala 27:21]
  assign FullAdder_82_io_b = io_B[82]; // @[Adder.scala 28:21]
  assign FullAdder_82_io_cin = FullAdder_81_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_83_io_a = io_A[83]; // @[Adder.scala 27:21]
  assign FullAdder_83_io_b = io_B[83]; // @[Adder.scala 28:21]
  assign FullAdder_83_io_cin = FullAdder_82_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_84_io_a = io_A[84]; // @[Adder.scala 27:21]
  assign FullAdder_84_io_b = io_B[84]; // @[Adder.scala 28:21]
  assign FullAdder_84_io_cin = FullAdder_83_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_85_io_a = io_A[85]; // @[Adder.scala 27:21]
  assign FullAdder_85_io_b = io_B[85]; // @[Adder.scala 28:21]
  assign FullAdder_85_io_cin = FullAdder_84_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_86_io_a = io_A[86]; // @[Adder.scala 27:21]
  assign FullAdder_86_io_b = io_B[86]; // @[Adder.scala 28:21]
  assign FullAdder_86_io_cin = FullAdder_85_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_87_io_a = io_A[87]; // @[Adder.scala 27:21]
  assign FullAdder_87_io_b = io_B[87]; // @[Adder.scala 28:21]
  assign FullAdder_87_io_cin = FullAdder_86_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_88_io_a = io_A[88]; // @[Adder.scala 27:21]
  assign FullAdder_88_io_b = io_B[88]; // @[Adder.scala 28:21]
  assign FullAdder_88_io_cin = FullAdder_87_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_89_io_a = io_A[89]; // @[Adder.scala 27:21]
  assign FullAdder_89_io_b = io_B[89]; // @[Adder.scala 28:21]
  assign FullAdder_89_io_cin = FullAdder_88_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_90_io_a = io_A[90]; // @[Adder.scala 27:21]
  assign FullAdder_90_io_b = io_B[90]; // @[Adder.scala 28:21]
  assign FullAdder_90_io_cin = FullAdder_89_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_91_io_a = io_A[91]; // @[Adder.scala 27:21]
  assign FullAdder_91_io_b = io_B[91]; // @[Adder.scala 28:21]
  assign FullAdder_91_io_cin = FullAdder_90_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_92_io_a = io_A[92]; // @[Adder.scala 27:21]
  assign FullAdder_92_io_b = io_B[92]; // @[Adder.scala 28:21]
  assign FullAdder_92_io_cin = FullAdder_91_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_93_io_a = io_A[93]; // @[Adder.scala 27:21]
  assign FullAdder_93_io_b = io_B[93]; // @[Adder.scala 28:21]
  assign FullAdder_93_io_cin = FullAdder_92_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_94_io_a = io_A[94]; // @[Adder.scala 27:21]
  assign FullAdder_94_io_b = io_B[94]; // @[Adder.scala 28:21]
  assign FullAdder_94_io_cin = FullAdder_93_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_95_io_a = io_A[95]; // @[Adder.scala 27:21]
  assign FullAdder_95_io_b = io_B[95]; // @[Adder.scala 28:21]
  assign FullAdder_95_io_cin = FullAdder_94_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_96_io_a = io_A[96]; // @[Adder.scala 27:21]
  assign FullAdder_96_io_b = io_B[96]; // @[Adder.scala 28:21]
  assign FullAdder_96_io_cin = FullAdder_95_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_97_io_a = io_A[97]; // @[Adder.scala 27:21]
  assign FullAdder_97_io_b = io_B[97]; // @[Adder.scala 28:21]
  assign FullAdder_97_io_cin = FullAdder_96_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_98_io_a = io_A[98]; // @[Adder.scala 27:21]
  assign FullAdder_98_io_b = io_B[98]; // @[Adder.scala 28:21]
  assign FullAdder_98_io_cin = FullAdder_97_io_cout; // @[Adder.scala 20:19 30:16]
  assign FullAdder_99_io_a = io_A[99]; // @[Adder.scala 27:21]
  assign FullAdder_99_io_b = io_B[99]; // @[Adder.scala 28:21]
  assign FullAdder_99_io_cin = FullAdder_98_io_cout; // @[Adder.scala 20:19 30:16]
endmodule
module Adder100(
  input         clock,
  input         reset,
  input  [99:0] a,
  input  [99:0] b,
  input         cin,
  output        cout,
  output [99:0] sum
);
  wire [99:0] myadder_io_A; // @[Adder100.scala 14:23]
  wire [99:0] myadder_io_B; // @[Adder100.scala 14:23]
  wire  myadder_io_Cin; // @[Adder100.scala 14:23]
  wire [99:0] myadder_io_Sum; // @[Adder100.scala 14:23]
  wire [99:0] myadder_io_Cout; // @[Adder100.scala 14:23]
  Adder myadder ( // @[Adder100.scala 14:23]
    .io_A(myadder_io_A),
    .io_B(myadder_io_B),
    .io_Cin(myadder_io_Cin),
    .io_Sum(myadder_io_Sum),
    .io_Cout(myadder_io_Cout)
  );
  assign cout = myadder_io_Cout[99]; // @[Adder100.scala 18:26]
  assign sum = myadder_io_Sum; // @[Adder100.scala 19:7]
  assign myadder_io_A = a; // @[Adder100.scala 15:16]
  assign myadder_io_B = b; // @[Adder100.scala 16:16]
  assign myadder_io_Cin = cin; // @[Adder100.scala 17:18]
endmodule
