module Q4i(
  output  out
);
  assign out = 1'h0; // @[Q4i.scala 8:7]
endmodule
