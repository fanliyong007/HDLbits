module MyWire(
  input   io_in,
  output  io_out
);
  assign io_out = io_in; // @[Wire.scala 39:10]
endmodule
